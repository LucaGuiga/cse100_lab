module hex7seg
    (input [3:0] N
    ,output [6:0] seg
    );

assign seg[0] = (~N[3] & ~N[2] & ~N[1] & N[0]) | (~N[3] & N[2] & ~N[1] & ~N[0]) | (N[3] & ~N[2] & N[1] & N[0]) | (N[3] & N[2] & ~N[1] & ~N[0]) | (N[3] & N[2] & ~N[1] & N[0]);
assign seg[1] = (~N[3] & ~N[2] & ~N[1] & N[0]) | (~N[3] & N[2] & ~N[1] & N[0]) | (~N[3] & N[2] & N[1] & ~N[0]) | (N[3] & ~N[2] & N[1] & N[0]) | (N[3] & N[2] & ~N[1] & ~N[0]) | (N[3] & N[2] & N[1] & ~N[0]) | (N[3] & N[2] & N[1] & N[0]);
assign seg[2] = (~N[3] & ~N[2] & ~N[1] & N[0]) | (~N[3] & ~N[2] & N[1] & ~N[0]) | (N[3] & N[2] & ~N[1] & ~N[0]) | (N[3] & N[2] & N[1] & ~N[0]) | (N[3] & N[2] & N[1] & N[0]);
assign seg[3] = (~N[3] & ~N[2] & ~N[1] & N[0]) | (~N[3] & N[2] & ~N[1] & ~N[0]) | (~N[3] & N[2] & N[1] & N[0]) | (N[3] & ~N[2] & ~N[1] & N[0]) | (N[3] & ~N[2] & N[1] & ~N[0]) | (N[3] & N[2] & N[1] & N[0]);
assign seg[4] = (~N[3] & ~N[2] & N[1] & N[0]) | (~N[3] & N[2] & ~N[1] & ~N[0]) | (~N[3] & N[2] & ~N[1] & N[0]) | (~N[3] & N[2] & N[1] & N[0]) | (N[3] & ~N[2] & ~N[1] & N[0]);
assign seg[5] = (~N[3] & ~N[2] & N[1] & ~N[0]) | (~N[3] & ~N[2] & N[1] & N[0]) | (~N[3] & N[2] & N[1] & N[0]) | (N[3] & N[2] & ~N[1] & ~N[0]) | (N[3] & N[2] & ~N[1] & N[0]);
assign seg[6] = (~N[3] & ~N[2] & ~N[1] & ~N[0]) | (~N[3] & ~N[2] & ~N[1] & N[0]);


endmodule


